`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    17:52:46 12/18/2020 
// Design Name: 
// Module Name:    Inst_Mem 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
`define BRANCH_TEST
module Inst_Mem(Address_in,Inst
    );
input [31:0] Address_in;
output wire[31:0] Inst;
reg [31:0] Rom[255:0];
assign Inst=Rom[Address_in[9:2]];
initial begin
`ifdef BASE_TEST
Rom[255]<=32'hffff_ffff;//idle instruction
Rom[0]<=32'b10001100000000010000000000000001; // Lw R1 1(R0)  
Rom[1]<=32'b10001100000000100000000000000010; // Lw R2 2(R0)  
Rom[2]<=32'b10001100000000110000000000000011; // Lw R3 3(R0)  
Rom[3]<=32'b10001100000001000000000000000100; // Lw R4 4(R0)  
Rom[4]<=32'b10001100000001010000000000000101; // Lw R5 5(R0)  
Rom[5]<=32'b00000000001000100010000000100000; // Add R4 R1 R2=>R4=R1+R2
Rom[6]<=32'b00000000001000110010100000100000; // Add R5 R1 R3=>R5=R1+R3
Rom[7]<=32'b10001100000000010000000000001010; // Lw R1 10(R0)  
Rom[8]<=32'b10001100001000100000000000000001; // Lw R2 1(R1) 
Rom[9]<=32'b10001100001000110000000000000010; // Lw R3 2(R1) 
Rom[10]<=32'b00000000011001000010100000100000; // Add R5 R3 R4=>R5=R3+R4
Rom[11]<=32'b00000000011000100011000000100000; // Add R6 R3 R2=>R6=R3+R2
Rom[12]<=32'b00000000110001110100100000100010; // Sub R9 R6 R7=>R9=R6-R7
Rom[13]<=32'b00000000110010000101000000100010; // Sub R10 R6 R8=>R10=R6-R8
Rom[14]<=32'b10001101010010110000000000000000; // Lw  R11 0(R10)
Rom[15]<=32'b10001101010011000000000000000010; // Lw  R12 2(R10)
`endif
`ifdef ADD_TEST_1
Rom[255]<=32'hffff_ffff;//idle instruction
Rom[0]<=32'b10001101011010100000000000000001; // Lw R10 1(R11) 
Rom[1]<=32'b10001101101011000000000000000001; // Lw R12 1(R13) 
Rom[2]<=32'b00000001100011000111000000100000; // Add R14 R12 R12=>R14=R12+R12

Rom[3]<=32'b10001101011010100000000000000010; // Lw R10 2(R11) 
Rom[4]<=32'b10001101101011000000000000000010; // Lw R12 2(R13) 
Rom[5]<=32'b00000001100010100111000000100000; // Add R14 R12 R10=>R14=R12+R10

Rom[6]<=32'b10001101011010100000000000000011; // Lw R10 3(R11) 
Rom[7]<=32'b10001101101011000000000000000011; // Lw R12 3(R13) 
Rom[8]<=32'b00000001010011000111000000100000; // Add R14 R10 R12=>R14=R10+R12

Rom[9]<=32'b10001101011010100000000000000100; // Lw R10 4(R11) 
Rom[10]<=32'b10001101101011000000000000000100; // Lw R12 4(R13) 
Rom[11]<=32'b00000001010010100111000000100000; // Add R14 R10 R10=>R14=R10+R10

Rom[12]<=32'b00000010000100010111100000100000; // Add R15 R16 R17=>R15=R16+R17
Rom[13]<=32'b00000010011101001001000000100000; // Add R18 R19 R20=>R18=R19+R20
Rom[14]<=32'b00000010010100100111100000100000; // Add R15 R18 R18=>R15=R18+R18

Rom[15]<=32'b00000010000100010111100000100000; // Add R15 R16 R17=>R15=R16+R17
Rom[16]<=32'b00000010011101001001000000100000; // Add R18 R19 R20=>R18=R19+R20
Rom[17]<=32'b00000010010011110111100000100000; // Add R15 R18 R15=>R15=R18+R15

Rom[18]<=32'b00000010000100010111100000100000; // Add R15 R16 R17=>R15=R16+R17
Rom[19]<=32'b00000010011101001001000000100000; // Add R18 R19 R20=>R18=R19+R20
Rom[20]<=32'b00000001111100101001000000100000; // Add R18 R15 R18=>R18=R15+R18

Rom[21]<=32'b00000010000100010111100000100000; // Add R15 R16 R17=>R15=R16+R17
Rom[22]<=32'b00000010011101001001000000100000; // Add R18 R19 R20=>R18=R19+R20
Rom[23]<=32'b00000001111011111001000000100000; // Add R18 R15 R15=>R18=R15+R15

`endif
`ifdef ADD_TEST_2
Rom[255]<=32'hffff_ffff;//idle instruction
Rom[0]<=32'b10001101011010100000000000000001; // Lw R10 1(R11) 
Rom[1]<=32'b00000001101011100110000000100000; // Add R12 R13 R14=>R12=R13+R14
Rom[2]<=32'b00000001100011000111100000100000; // Add R15 R12 R12=>R15=R12+R12

Rom[3]<=32'b10001101011010100000000000000010; // Lw R10 2(R11) 
Rom[4]<=32'b00000001101011100110000000100000; // Add R12 R13 R14=>R12=R13+R14
Rom[5]<=32'b00000001100010100111100000100000; // Add R15 R12 R10=>R15=R12+R10

Rom[6]<=32'b10001101011010100000000000000011; // Lw R10 3(R11) 
Rom[7]<=32'b00000001101011100110000000100000; // Add R12 R13 R14=>R12=R13+R14
Rom[8]<=32'b00000001010011000111100000100000; // Add R15 R10 R12=>R15=R10+R12

Rom[9]<=32'b10001101011010100000000000000100; // Lw R10 4(R11) 
Rom[10]<=32'b00000001101011100110000000100000; // Add R12 R13 R14=>R12=R13+R14
Rom[11]<=32'b00000001010010100111100000100000; // Add R15 R10 R10=>R15=R10+R10

Rom[12]<=32'b00000010001100101000000000100000; // Add R16 R17 R18=>R16=R17+R18
Rom[13]<=32'b10001110100100110000000000000001; // Lw R19 1(R20) 
Rom[14]<=32'b00000010011100110101000000100000; // Add R10 R19 R19=>R10=R19+R19

Rom[15]<=32'b00000010001100101000000000100000; // Add R16 R17 R18=>R16=R17+R18
Rom[16]<=32'b10001110100100110000000000000010; // Lw R19 2(R20) 
Rom[17]<=32'b00000010011100000101000000100000; // Add R10 R19 R16=>R10=R19+R16

Rom[18]<=32'b00000010001100101000000000100000; // Add R16 R17 R18=>R16=R17+R18
Rom[19]<=32'b10001110100100110000000000000011; // Lw R19 3(R20) 
Rom[20]<=32'b00000010000100110101000000100000; // Add R10 R16 R19=>R10=R16+R19

Rom[21]<=32'b00000010001100101000000000100000; // Add R16 R17 R18=>R16=R17+R18
Rom[22]<=32'b10001110100100110000000000000100; // Lw R19 4(R20) 
Rom[23]<=32'b00000010000100000101000000100000; // Add R10 R16 R16=>R10=R16+R16
`endif
`ifdef BRANCH_TEST  //R5 is i ,R1 is j
Rom[255]<=32'hffff_ffff;//idle instruction
Rom[0]<=32'b00000000101000100010100000100000;  //Add R5 R5 R2
Rom[1]<=32'b00000000001000010000100000100010; // Sub R1 R1 R1=>R1=0
Rom[2]<=32'b00000000001000100000100000100000;  //Add R1 R1 R2
Rom[3]<=32'b00000000100000010001100000101010; // slt R3 R4 R1=>R3=R4<=R1?1:0
Rom[4]<=32'hffff_ffff;
Rom[5]<=32'b00010000000000111111111111111101; // beq R0 R3 -3
Rom[6]<=32'b00000000110001010011100000101010; // slt R7 R6 R5=>R7=R6<=R5?1:0
Rom[7]<=32'hffff_ffff;
Rom[8]<=32'b00010000000001111111111111111000; // beq R0 R7 -8
`endif
end
endmodule
